module DIV(
	Y,
	A,
	B,
	aDiv
);

output wire [7:0] Y;
input wire [3:0] A;
input wire [3:0] B;
input wire aDiv;

endmodule
